LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_unsigned.ALL;

ENTITY LED_7SEG IS
	GENERIC(
		DATA_LENGTH	: INTEGER
	);
	PORT(
		I_CLK 	: IN 	STD_LOGIC;
		I_DATA	: IN  STD_LOGIC_VECTOR(DATA_LENGTH - 1 DOWNTO 0);
		O_LED7	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEHAVIORAL OF LED_7SEG IS

BEGIN
	PROCESS(I_CLK)
	BEGIN
		IF (I_DATA = "0000") THEN-------0
			O_LED7 <= "11000000";
		ELSIF(I_DATA = "0001") THEN-----1
			O_LED7 <= "11111001";
		ELSIF(I_DATA = "0010") THEN-----2
			O_LED7 <= "10100100";
		ELSIF(I_DATA = "0011") THEN-----3
			O_LED7 <= "10110000";
		ELSIF(I_DATA = "0100") THEN-----4
			O_LED7 <= "10011001";
		ELSIF(I_DATA = "0101") THEN-----5
			O_LED7 <= "10010010";
		ELSIF(I_DATA = "0110") THEN-----6
			O_LED7 <= "10000010";
		ELSIF(I_DATA = "0111") THEN-----7
			O_LED7 <= "11111000";
		ELSIF(I_DATA = "1000") THEN-----8
			O_LED7 <= "10000000";
		ELSIF(I_DATA = "1001") THEN-----9
			O_LED7 <= "10010000";
		END IF; 
	END PROCESS;
END ARCHITECTURE;
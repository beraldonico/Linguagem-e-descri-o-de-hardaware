LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY CAMINHO_DADOS IS
	GENERIC(
		P_DATA	: INTEGER	:= 8
	);
	PORT(
		I_CLK			:  IN STD_LOGIC;
		I_RST			:  IN STD_LOGIC;
		I_WE			:  IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		I_DATA		:  IN STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0);
		I_SEL_RS1	:  IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		I_SEL_RS2	:  IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		I_SEL_ULA	:  IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		I_SEL_IMED	:	IN STD_LOGIC;
		I_EN_OUT		:	IN STD_LOGIC;
		O_LED			: OUT STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEHAVIORAL OF CAMINHO_DADOS IS
	COMPONENT BANCO_DE_REGISTRADORES IS
		GENERIC(
			P_DATA	: INTEGER := 8
		);
		PORT(
			I_CLK			:  IN STD_LOGIC;
			I_RST			:  IN STD_LOGIC;
			I_WE			:  IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			I_DATA		:  IN STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0);
			I_SEL_RS1	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			I_SEL_RS2	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			O_RS1			: OUT STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0);
			O_RS2			: OUT STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0)
		);
	END COMPONENT;
	
	COMPONENT ULA IS
		GENERIC(
			P_DATA	:	INTEGER := 16
		);
		PORT(
			I_SEL	:  IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			I_RS1	:  IN STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0);
			I_RS2	:  IN STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0);
			O_ULA	: OUT STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0)
		);
	END COMPONENT;
	
	SIGNAL W_RS1	: STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0);
	SIGNAL W_RS2	: STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0);
	SIGNAL W_ULA	: STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0);
	SIGNAL W_DATA	: STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0);
	
	COMPONENT REGISTRADOR IS
		GENERIC(
			P_DATA	: INTEGER := 16
		);
		PORT(
			I_CLK		:  IN STD_LOGIC;
			I_RST		:  IN STD_LOGIC;
			I_WE		:  IN STD_LOGIC;
			I_DATA	:  IN STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0);
			O_DATA	: OUT STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0) 
		);
	END COMPONENT;
	
BEGIN
	
	W_DATA <= I_DATA WHEN (I_SEL_IMED = '0') ELSE W_ULA;

	U00 : BANCO_DE_REGISTRADORES
		GENERIC MAP(
      	P_DATA	=> P_DATA
      )
		PORT MAP(
      	I_CLK			=> I_CLK,
      	I_RST			=> I_RST,
      	I_WE			=> I_WE,
      	I_DATA		=> W_DATA,
      	I_SEL_RS1	=> I_SEL_RS1,
      	I_SEL_RS2	=> I_SEL_RS2,
      	O_RS1			=> W_RS1,
      	O_RS2			=> W_RS2
		);
		
	U01 : ULA
		GENERIC MAP(
			P_DATA => P_DATA
		)
		PORT MAP(
			I_SEL	=> I_SEL_ULA,
			I_RS1	=> W_RS1,
			I_RS2	=> W_RS2,
			O_ULA	=> W_ULA
		); 
		
	U02 : REGISTRADOR
		GENERIC MAP(
			P_DATA	=> P_DATA
		)
		PORT MAP(
			I_CLK		=> I_CLK, 
			I_RST		=> I_RST,
			I_WE		=> I_EN_OUT,
			I_DATA	=> W_ULA,
			O_DATA	=> O_LED
		);
END ARCHITECTURE;
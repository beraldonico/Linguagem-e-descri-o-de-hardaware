LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_unsigned.ALL;

ENTITY MEMORIA IS
	GENERIC(
		DATA_LENGTH	: INTEGER;
		ADD_LENGTH	: INTEGER
	);
	PORT(
		I_CLK 	: IN 	STD_LOGIC;
		I_WE		: IN  STD_LOGIC;
		I_ADD 	: IN  STD_LOGIC_VECTOR(ADD_LENGTH - 1 DOWNTO 0);
		I_DATA	: IN  STD_LOGIC_VECTOR(DATA_LENGTH - 1 DOWNTO 0);
		O_DATA	: OUT STD_LOGIC_VECTOR(DATA_LENGTH - 1 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEHAVIORAL OF MEMORIA IS
	TYPE MEM_TYPE IS ARRAY(2**ADD_LENGTH-1 DOWNTO 0) OF STD_LOGIC_VECTOR(DATA_LENGTH-1 DOWNTO 0);
	SIGNAL W_MEMORIA_RAM : MEM_TYPE;
BEGIN
	PROCESS(I_CLK)
	BEGIN
		IF(I_WE = '1')THEN
			W_MEMORIA_RAM(CONV_INTEGER(I_ADD)) <= I_DATA;
		ELSE
			O_DATA <= W_MEMORIA_RAM(CONV_INTEGER(I_ADD));
		END IF;
	END PROCESS;
END ARCHITECTURE;
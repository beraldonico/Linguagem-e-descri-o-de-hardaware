LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FLIP_FLOP_32 IS
	GENERIC(
		S_DATA  : INTEGER := 32
	);
	PORT(
		I_DATA  : IN  STD_LOGIC_VECTOR(S_DATA - 1 DOWNTO 0);
		I_RST   : IN  STD_LOGIC;
		I_EN    : IN  STD_LOGIC;
		I_CLK   : IN  STD_LOGIC;
		O_DATA  : OUT STD_LOGIC_VECTOR(S_DATA - 1 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEHAVIORAL OF FLIP_FLOP_32 IS

BEGIN
	PROCESS(I_CLK, I_RST)
		BEGIN
			IF (I_EN = '1') THEN
				IF (I_RST = '1') THEN
					O_DATA <= (OTHERS => '0');
				ELSIF RISING_EDGE(I_CLK) THEN
					O_DATA <= I_DATA;
				END IF;
			END IF;
		END PROCESS;
END ARCHITECTURE;
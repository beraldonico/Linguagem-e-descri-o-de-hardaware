LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_unsigned.ALL;

ENTITY STMEMORIA IS
	PORT(
		I_CLK		: IN  STD_LOGIC;
		I_BTNW	: IN  STD_LOGIC;
		I_BTNR	: IN  STD_LOGIC;
		I_BTNRST	: IN  STD_LOGIC;
		O_WE		: OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE BEHAVIORAL OF STMEMORIA IS
	TYPE STATE_TYPE IS (ST_IDLE, ST_WRITE, ST_READ);
	SIGNAL STATE : STATE_TYPE := ST_IDLE;
BEGIN
	PROCESS(I_CLK, I_BTNRST)
	BEGIN
		IF(I_BTNRST = '0') THEN
				O_WE <= '0';
				STATE <= ST_IDLE;
				--o que falta
		ELSIF RISING_EDGE (I_CLK) THEN
			CASE STATE IS
				WHEN ST_IDLE =>
					IF(I_BTNR = '0')THEN
						O_WE <= '0';
						STATE <= ST_READ;
					ELSIF(I_BTNW = '0')THEN
						O_WE <= '1';
						STATE <= ST_WRITE;
					ELSE
						O_WE <= '0';
						STATE <= ST_IDLE;
					END IF;
				WHEN ST_READ =>
					IF(I_BTNR = '1')THEN
						O_WE <= '0';
						STATE <= ST_IDLE;
					END IF;
				WHEN ST_WRITE =>
					IF(I_BTNW = '1')THEN
						O_WE <= '0';
						STATE <= ST_IDLE;
					END IF;
				WHEN OTHERS =>
					NULL;
			END CASE;
		END IF;
	END PROCESS;
END ARCHITECTURE;
--TB_TRABALHO_STMEMORIA/TBTSTM/W_WE		|NO DATA ?!?!?!?!?!?
--TB_TRABALHO_STMEMORIA/TBTSTM/W_DATA	|
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_unsigned.ALL;

ENTITY TRABALHO_STMEMORIA IS
	GENERIC(
		DATA_LENGTH	: INTEGER := 4;
		ADD_LENGTH	: INTEGER := 5
	);
	PORT(
		I_CLK		: IN  STD_LOGIC;
		I_BTNW	: IN  STD_LOGIC;
		I_BTNR	: IN  STD_LOGIC;
		I_BTNRST	: IN  STD_LOGIC;
		I_ADD 	: IN  STD_LOGIC_VECTOR(ADD_LENGTH - 1 DOWNTO 0);
		I_DATA	: IN  STD_LOGIC_VECTOR(DATA_LENGTH - 1 DOWNTO 0);
		O_LED7	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEHAVIORAL OF TRABALHO_STMEMORIA IS
	COMPONENT STMEMORIA IS
		PORT(
		I_CLK		: IN  STD_LOGIC;
		I_BTNW	: IN  STD_LOGIC;
		I_BTNR	: IN  STD_LOGIC;
		I_BTNRST	: IN  STD_LOGIC;
		O_WE		: OUT STD_LOGIC
	);
	END COMPONENT;
	SIGNAL W_WE	: STD_LOGIC;
	
	COMPONENT MEMORIA IS
		GENERIC(
			DATA_LENGTH	: INTEGER;
			ADD_LENGTH	: INTEGER
		);
		PORT(
			I_CLK 	: IN 	STD_LOGIC;
			I_WE		: IN  STD_LOGIC;
			I_ADD 	: IN  STD_LOGIC_VECTOR(ADD_LENGTH - 1 DOWNTO 0);
			I_DATA	: IN  STD_LOGIC_VECTOR(DATA_LENGTH - 1 DOWNTO 0);
			O_DATA	: OUT STD_LOGIC_VECTOR(DATA_LENGTH - 1 DOWNTO 0)
		);
	END COMPONENT;
	SIGNAL W_DATA : STD_LOGIC_VECTOR(DATA_LENGTH - 1 DOWNTO 0);
	
	COMPONENT LED_7SEG IS
		GENERIC(
			DATA_LENGTH	: INTEGER
		);
		PORT(
			I_CLK 	: IN 	STD_LOGIC;
			I_DATA	: IN  STD_LOGIC_VECTOR(DATA_LENGTH - 1 DOWNTO 0);
			O_LED7	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
	END COMPONENT;
	
BEGIN
	ST : STMEMORIA
		PORT MAP(
			I_CLK			=> I_CLK,
			I_BTNW		=> I_BTNR,
			I_BTNR		=> I_BTNW,
			I_BTNRST		=> I_BTNRST,
			O_WE			=> W_WE
		);	
	RAM : MEMORIA
		GENERIC MAP(
			DATA_LENGTH => DATA_LENGTH,
			ADD_LENGTH	=> ADD_LENGTH
		)
		PORT MAP(
			I_CLK  => I_CLK,
			I_WE 	 => W_WE,
			I_ADD  => I_ADD,
			I_DATA => I_DATA,
			O_DATA => W_DATA
		);
	LED : LED_7SEG
		GENERIC MAP(
			DATA_LENGTH => DATA_LENGTH
		)
		PORT MAP(
			I_CLK	 => I_CLK,
			I_DATA => W_DATA,
			O_LED7 => O_LED7
		);
END ARCHITECTURE;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY BANCO_DE_REGISTRADORES IS
	GENERIC(
		P_DATA	: INTEGER := 8
	);
	PORT(
		I_CLK			:  IN STD_LOGIC;
		I_RST			:  IN STD_LOGIC;
		I_WE			:  IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		I_DATA		:  IN STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0);
		I_SEL_RS1	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		I_SEL_RS2	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		O_RS1			: OUT STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0);
		O_RS2			: OUT STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEHAVIORAL OF BANCO_DE_REGISTRADORES IS
	COMPONENT REGISTRADOR IS
		GENERIC(
			P_DATA	: INTEGER := 16
		);
		PORT(
			I_CLK		:  IN STD_LOGIC;
			I_RST		:  IN STD_LOGIC;
			I_WE		:  IN STD_LOGIC;
			I_DATA	:  IN STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0);
			O_DATA	: OUT STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0) 
		);
	END COMPONENT;
	COMPONENT MULTIPLEXADOR IS
		GENERIC(
			P_DATA	: INTEGER := 16
		);
		
		PORT(
			I_SEL  	:	 IN STD_LOGIC_VECTOR(1 downto 0);
			I_DATA0	:	 IN STD_LOGIC_VECTOR(p_DATA-1 downto 0);
			I_DATA1	:	 IN STD_LOGIC_VECTOR(p_DATA-1 downto 0);
			I_DATA2	:	 IN STD_LOGIC_VECTOR(p_DATA-1 downto 0);
			I_DATA3	:	 IN STD_LOGIC_VECTOR(p_DATA-1 downto 0);
			O_DATA 	:	OUT STD_LOGIC_VECTOR(p_DATA-1 downto 0)
			
		);
	END COMPONENT;
	
	SIGNAL W_DATA0	:	STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0);
	SIGNAL W_DATA1	:	STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0);
	SIGNAL W_DATA2	:	STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0);
	SIGNAL W_DATA3	:	STD_LOGIC_VECTOR(P_DATA - 1 DOWNTO 0);
	
BEGIN
	
	UR0 : REGISTRADOR
		GENERIC MAP(
			P_DATA => P_DATA
		)
		PORT MAP(
			I_CLK	 => I_CLK,
			I_RST	 => I_RST,
			I_WE	 => I_WE(0),
			I_DATA => I_DATA,
		   O_DATA => W_DATA0
		);
	UR1 : REGISTRADOR
		GENERIC MAP(
			P_DATA => P_DATA
		)
		PORT MAP(
			I_CLK	 => I_CLK,
			I_RST	 => I_RST,
			I_WE	 => I_WE(1),
			I_DATA => I_DATA,
		   O_DATA => W_DATA1
		);
	UR2 : REGISTRADOR
		GENERIC MAP(
			P_DATA => P_DATA
		)
		PORT MAP(
			I_CLK	 => I_CLK,
			I_RST	 => I_RST,
			I_WE	 => I_WE(2),
			I_DATA => I_DATA,
		   O_DATA => W_DATA2
		);
	UR3 : REGISTRADOR
		GENERIC MAP(
			P_DATA => P_DATA
		)
		PORT MAP(
			I_CLK	 => I_CLK,
			I_RST	 => I_RST,
			I_WE	 => I_WE(3),
			I_DATA => I_DATA,
		   O_DATA => W_DATA3
		);
		
	MUX1 : MULTIPLEXADOR
		GENERIC MAP(
			P_DATA	=> P_DATA
		)
		PORT MAP(
			I_SEL  	=> I_SEL_RS1,
			I_DATA0	=> W_DATA0,
			I_DATA1	=> W_DATA1,
			I_DATA2	=> W_DATA2,
			I_DATA3	=> W_DATA3,
			O_DATA 	=> O_RS1
			
		);
		
	MUX2 : MULTIPLEXADOR
		GENERIC MAP(
			P_DATA	=> P_DATA
		)
		PORT MAP(
			I_SEL  	=> I_SEL_RS2,
			I_DATA0	=> W_DATA0,
			I_DATA1	=> W_DATA1,
			I_DATA2	=> W_DATA2,
			I_DATA3	=> W_DATA3,
			O_DATA 	=> O_RS2
			
		);	
	
END ARCHITECTURE;